class array_bfm;
	
endclass

