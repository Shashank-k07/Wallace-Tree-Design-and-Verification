class axi_tx;
	randc bit[3:0]a,b;
endclass
